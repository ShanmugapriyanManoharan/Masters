library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package arraypackage is
type Memory_Array is array (0 to 29) of STD_LOGIC_VECTOR (31 downto 0);
end arraypackage;